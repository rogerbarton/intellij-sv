timeunit 1us;
timeprecision 1ps;

module empty ();

endmodule

extern module ext1;

module empty2 #() ();

endmodule

extern module ext2 #() ();

module empty3 #(
    parameter unsigned Order
) ();

endmodule

module empty3 #() (
    input logic clk_i
);

endmodule


module empty3 #(
    parameter unsigned Order
) (
    input logic clk_i
);

endmodule


module filter #(
//    parameter int unsigned Order      = 127, // Filter order
//    parameter int unsigned AddrWidth  = 7   // Address width
  ) (
    input logic clk_i,                         // Clock signal

    input logic                 data_in_req_i, // Req at input
    input logic [DataWidth-1:0] data_in_i,     // Incoming data
  );

endmodule : filter