timeunit 1us;
timeunit
timeunit 1s;
timeunit ;
timeunit 1us/;
timeunit 0s/9ps;
timeprecision 1ps;
